package struct_define;
    
endpackage
